module reciep_MLUT (
    input logic [3:0] selector,
    output logic [15:0] value
);

always_comb 
begin  
    case(selector)
        // 'd0: value = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        // 'd1: value = 64'b1111111110000000000000000000000000000000000000000000000000000000;
        // 'd2: value = 64'b1111111111010101010101010101010101000111000001000100101101101010;
        // 'd3: value = 64'b1111111111101010101010101010101010111000111110111011010010010111;
        // 'd4: value = 64'b1111111111110011001100110011001100110011001100110011001100110011;
         
        'd0: value = 16'b1000000001000001;
        'd1: value = 16'b1111111111100000;
        'd2: value = 16'b1111111111110110;
        'd3: value = 16'b1111111111111011;
        'd4: value = 16'b1111111111111101;

        'd5: value = 16'b1111111111111110;
        'd6: value = 16'b1111111111111111;
        'd7: value = 16'b1111111111111111;
        'd8: value = 16'b0;
        'd9: value = 16'b0; 
              
        default:
        value = 'b0;
         
    endcase
    
end


endmodule


module reciep_CLUT (
    input logic [3:0] selector,
    output logic [31:0] value
);

always_comb 
begin  
    case(selector)
        // 'd0: value = 64'b0111111111111111000000000000000000000000000000000000000000000000;
        // 'd1: value = 64'b0000000001100000000000000000000000000000000000000000000000000000;
        // 'd2: value = 64'b0000000000110101010101010101010101010001110000010001001011011010;
        // 'd3: value = 64'b0000000000100101010101010101010101010001110000010001001011011010;
        // 'd4: value = 64'b0000000000011100110011001100110011001100110011001100110011001101;

        'd0: value = 32'b00000000000111111111111111000000;
        'd1: value = 32'b00000000000000000001100000000000;
        'd2: value = 32'b00000000000000000000110101010101;
        'd3: value = 32'b00000000000000000000100101010101;
        'd4: value = 32'b00000000000000000000011100110011;

        'd5: value = 32'b00000000000000000000010111011101;
        'd6: value = 32'b00000000000000000000010001001001;
        'd7: value = 32'b00000000000000000000110101010101;
        'd8: value = 32'b00000000000000000000001111000111;
        'd9: value = 32'b00000000000000000000001101100000;
        default:
        value = 'b0;
         
    endcase
    
end


endmodule